module my_or (output out, input in1, in2);

	or or1(out, in1, in2);

endmodule