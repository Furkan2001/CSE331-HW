module my_xor_32_bit (output [31:0] out, input [31:0] in1, in2);

	my_xor xor1 (out[0], in1[0], in2[0]);
	my_xor xor2 (out[1], in1[1], in2[1]);
	my_xor xor3 (out[2], in1[2], in2[2]);
	my_xor xor4 (out[3], in1[3], in2[3]);
	my_xor xor5 (out[4], in1[4], in2[4]);
	my_xor xor6 (out[5], in1[5], in2[5]);
	my_xor xor7 (out[6], in1[6], in2[6]);
	my_xor xor8 (out[7], in1[7], in2[7]);
	my_xor xor9 (out[8], in1[8], in2[8]);
	my_xor xor10 (out[9], in1[9], in2[9]);
	my_xor xor11 (out[10], in1[10], in2[10]);
	my_xor xor12 (out[11], in1[11], in2[11]);
	my_xor xor13 (out[12], in1[12], in2[12]);
	my_xor xor14 (out[13], in1[13], in2[13]);
	my_xor xor15 (out[14], in1[14], in2[14]);
	my_xor xor16 (out[15], in1[15], in2[15]);
	my_xor xor17 (out[16], in1[16], in2[16]);
	my_xor xor18 (out[17], in1[17], in2[17]);
	my_xor xor19 (out[18], in1[18], in2[18]);
	my_xor xor20 (out[19], in1[19], in2[19]);
	my_xor xor21 (out[20], in1[20], in2[20]);
	my_xor xor22 (out[21], in1[21], in2[21]);
	my_xor xor23 (out[22], in1[22], in2[22]);
	my_xor xor24 (out[23], in1[23], in2[23]);
	my_xor xor25 (out[24], in1[24], in2[24]);
	my_xor xor26 (out[25], in1[25], in2[25]);
	my_xor xor27 (out[26], in1[26], in2[26]);
	my_xor xor28 (out[27], in1[27], in2[27]);
	my_xor xor29 (out[28], in1[28], in2[28]);
	my_xor xor30 (out[29], in1[29], in2[29]);
	my_xor xor31 (out[30], in1[30], in2[30]);
	my_xor xor32 (out[31], in1[31], in2[31]);

endmodule