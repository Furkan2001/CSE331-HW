module design_p_and_g (output [31:0] G1, P1, output [7:0] G2, P2, input [31:0] A, B);
	wire x0,x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23;

	and and1(G1[0], A[0], B[0]);
	or or1(P1[0], A[0], B[0]);

	and and2(G1[1], A[1], B[1]);
	or or2(P1[1], A[1], B[1]);

	and and3(G1[2], A[2], B[2]);
	or or3(P1[2], A[2], B[2]);

	and and4(G1[3], A[3], B[3]);
	or or4(P1[3], A[3], B[3]);

	// G3:0 = g3 + p3g2 + p3p2g1 + p3p2p1g0
	// P3:0 = p3p2p1p0
	and and33(x0, G1[0], P1[1], P1[2], P1[3]); 
	and and34(x1, P1[3], P1[2], G1[1]);
	and and35(x2, P1[3], G1[2]);
	or or33(G2[0], G1[3], x0, x1, x2); //G3:0
	and and36(P2[0], P1[0], P1[1], P1[2], P1[3]); //P3:0

	and and5(G1[4], A[4], B[4]);
	or or5(P1[4], A[4], B[4]);

	and and6(G1[5], A[5], B[5]);
	or or6(P1[5], A[5], B[5]);

	and and7(G1[6], A[6], B[6]);
	or or7(P1[6], A[6], B[6]);

	and and8(G1[7], A[7], B[7]);
	or or8(P1[7], A[7], B[7]);

	and and37(x3, G1[4], P1[5], P1[6], P1[7]); 
	and and38(x4, P1[7], P1[6], G1[5]);
	and and39(x5, P1[7], G1[6]);
	or or34(G2[1], G1[7], x3, x4, x5); //G7:4
	and and40(P2[1], P1[4], P1[5], P1[6], P1[7]); //P7:4

	and and9(G1[8], A[8], B[8]);
	or or9(P1[8], A[8], B[8]);

	and and10(G1[9], A[9], B[9]);
	or or10(P1[9], A[9], B[9]);

	and and11(G1[10], A[10], B[10]);
	or or11(P1[10], A[10], B[10]);

	and and12(G1[11], A[11], B[11]);
	or or12(P1[11], A[11], B[11]);

	and and41(x6, G1[8], P1[9], P1[10], P1[11]); 
	and and42(x7, P1[11], P1[10], G1[9]);
	and and43(x8, P1[11], G1[10]);
	or or35(G2[2], G1[11], x6, x7, x8); //G11:8
	and and44(P2[2], P1[8], P1[9], P1[10], P1[11]); //P11:8

	and and13(G1[12], A[12], B[12]);
	or or13(P1[12], A[12], B[12]);

	and and14(G1[13], A[13], B[13]);
	or or14(P1[13], A[13], B[13]);

	and and15(G1[14], A[14], B[14]);
	or or15(P1[14], A[14], B[14]);

	and and16(G1[15], A[15], B[15]);
	or or16(P1[15], A[15], B[15]);

	and and45(x9, G1[12], P1[13], P1[14], P1[15]); 
	and and46(x10, P1[15], P1[14], G1[13]);
	and and47(x11, P1[15], G1[14]);
	or or36(G2[3], G1[15], x9, x10, x11); //G15:12
	and and48(P2[3], P1[12], P1[13], P1[14], P1[15]); //P15:12

	and and17(G1[16], A[16], B[16]);
	or or17(P1[16], A[16], B[16]);

	and and18(G1[17], A[17], B[17]);
	or or18(P1[17], A[17], B[17]);

	and and19(G1[18], A[18], B[18]);
	or or19(P1[18], A[18], B[18]);

	and and20(G1[19], A[19], B[19]);
	or or20(P1[19], A[19], B[19]);

	and and49(x12, G1[16], P1[17], P1[18], P1[19]); 
	and and50(x13, P1[19], P1[18], G1[17]);
	and and51(x14, P1[19], G1[18]);
	or or37(G2[4], G1[19], x12, x13, x14); //G19:16
	and and52(P2[4], P1[16], P1[17], P1[18], P1[19]); //P19:16

	and and21(G1[20], A[20], B[20]);
	or or21(P1[20], A[20], B[20]);

	and and22(G1[21], A[21], B[21]);
	or or22(P1[21], A[21], B[21]);

	and and23(G1[22], A[22], B[22]);
	or or23(P1[22], A[22], B[22]);

	and and24(G1[23], A[23], B[23]);
	or or24(P1[23], A[23], B[23]);

	and and53(x15, G1[20], P1[21], P1[22], P1[23]); 
	and and54(x16, P1[23], P1[22], G1[21]);
	and and55(x17, P1[23], G1[22]);
	or or38(G2[5], G1[23], x15, x16, x17); //G23:20
	and and56(P2[5], P1[20], P1[21], P1[22], P1[23]); //P23:20

	and and25(G1[24], A[24], B[24]);
	or or25(P1[24], A[24], B[24]);

	and and26(G1[25], A[25], B[25]);
	or or26(P1[25], A[25], B[25]);

	and and27(G1[26], A[26], B[26]);
	or or27(P1[26], A[26], B[26]);

	and and28(G1[27], A[27], B[27]);
	or or28(P1[27], A[27], B[27]);

	and and57(x18, G1[24], P1[25], P1[26], P1[27]); 
	and and58(x19, P1[27], P1[26], G1[25]);
	and and59(x20, P1[27], G1[26]);
	or or39(G2[6], G1[27], x18, x19, x20); //G27:24
	and and60(P2[6], P1[24], P1[25], P1[26], P1[27]); //P27:24

	and and29(G1[28], A[28], B[28]);
	or or29(P1[28], A[28], B[28]);

	and and30(G1[29], A[29], B[29]);
	or or30(P1[29], A[29], B[29]);

	and and31(G1[30], A[30], B[30]);
	or or31(P1[30], A[30], B[30]);

	and and32(G1[31], A[31], B[31]);
	or or32(P1[31], A[31], B[31]);

	and and61(x21, G1[28], P1[29], P1[30], P1[31]); 
	and and62(x22, P1[31], P1[30], G1[29]);
	and and63(x23, P1[31], G1[30]);
	or or40(G2[7], G1[31], x21, x22, x23); //G31:28
	and and64(P2[7], P1[28], P1[29], P1[30], P1[31]); //P31:28

 

endmodule
