module my_and (output out, input in1, in2);

	and and1(out, in1, in2);

endmodule
