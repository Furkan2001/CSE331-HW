module my_xor (output out, input in1, in2);

	xor xor1(out, in1, in2);

endmodule